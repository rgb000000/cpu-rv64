module SimTop(
  input         clock,
  input         reset,
  input  [63:0] io_logCtrl_log_begin,
  input  [63:0] io_logCtrl_log_end,
  input  [63:0] io_logCtrl_log_level,
  input         io_perfInfo_clean,
  input         io_perfInfo_dump,
  output        io_uart_out_valid,
  output [7:0]  io_uart_out_ch,
  output        io_uart_in_valid,
  input  [7:0]  io_uart_in_ch,
  input         io_memAXI_0_aw_ready,
  output        io_memAXI_0_aw_valid,
  output [63:0] io_memAXI_0_aw_bits_addr,
  output [2:0]  io_memAXI_0_aw_bits_prot,
  output [3:0]  io_memAXI_0_aw_bits_id,
  output        io_memAXI_0_aw_bits_user,
  output [7:0]  io_memAXI_0_aw_bits_len,
  output [2:0]  io_memAXI_0_aw_bits_size,
  output [1:0]  io_memAXI_0_aw_bits_burst,
  output        io_memAXI_0_aw_bits_lock,
  output [3:0]  io_memAXI_0_aw_bits_cache,
  output [3:0]  io_memAXI_0_aw_bits_qos,
  input         io_memAXI_0_w_ready,
  output        io_memAXI_0_w_valid,
  output [63:0] io_memAXI_0_w_bits_data [3: 0],
  output [7:0]  io_memAXI_0_w_bits_strb,
  output        io_memAXI_0_w_bits_last,
  output        io_memAXI_0_b_ready,
  input         io_memAXI_0_b_valid,
  input  [1:0]  io_memAXI_0_b_bits_resp,
  input  [3:0]  io_memAXI_0_b_bits_id,
  input         io_memAXI_0_b_bits_user,
  input         io_memAXI_0_ar_ready,
  output        io_memAXI_0_ar_valid,
  output [63:0] io_memAXI_0_ar_bits_addr,
  output [2:0]  io_memAXI_0_ar_bits_prot,
  output [3:0]  io_memAXI_0_ar_bits_id,
  output        io_memAXI_0_ar_bits_user,
  output [7:0]  io_memAXI_0_ar_bits_len,
  output [2:0]  io_memAXI_0_ar_bits_size,
  output [1:0]  io_memAXI_0_ar_bits_burst,
  output        io_memAXI_0_ar_bits_lock,
  output [3:0]  io_memAXI_0_ar_bits_cache,
  output [3:0]  io_memAXI_0_ar_bits_qos,
  output        io_memAXI_0_r_ready,
  input         io_memAXI_0_r_valid,
  input  [1:0]  io_memAXI_0_r_bits_resp,
  input  [63:0] io_memAXI_0_r_bits_data [3: 0],
  input         io_memAXI_0_r_bits_last,
  input  [3:0]  io_memAXI_0_r_bits_id,
  input         io_memAXI_0_r_bits_user
);
  MySimTop mysimtop(
    .clock(clock),
    .reset(reset),
    .io_logCtrl_log_begin(io_logCtrl_log_begin),
    .io_logCtrl_log_end(io_logCtrl_log_end),
    .io_logCtrl_log_level(io_logCtrl_log_level),
    .io_perfInfo_clean(io_perfInfo_clean),
    .io_perfInfo_dump(io_perfInfo_dump),
    .io_uart_out_valid(io_uart_out_valid),
    .io_uart_out_ch(io_uart_out_ch),
    .io_uart_in_valid(io_uart_in_valid),
    .io_uart_in_ch(io_uart_in_ch),
    .io_memAXI_0_aw_ready(io_memAXI_0_aw_ready),
    .io_memAXI_0_aw_valid(io_memAXI_0_aw_valid),
    .io_memAXI_0_aw_bits_addr(io_memAXI_0_aw_bits_addr),
    .io_memAXI_0_aw_bits_prot(io_memAXI_0_aw_bits_prot),
    .io_memAXI_0_aw_bits_id(io_memAXI_0_aw_bits_id),
    .io_memAXI_0_aw_bits_user(io_memAXI_0_aw_bits_user),
    .io_memAXI_0_aw_bits_len(io_memAXI_0_aw_bits_len),
    .io_memAXI_0_aw_bits_size(io_memAXI_0_aw_bits_size),
    .io_memAXI_0_aw_bits_burst(io_memAXI_0_aw_bits_burst),
    .io_memAXI_0_aw_bits_lock(io_memAXI_0_aw_bits_lock),
    .io_memAXI_0_aw_bits_cache(io_memAXI_0_aw_bits_cache),
    .io_memAXI_0_aw_bits_qos(io_memAXI_0_aw_bits_qos),
    .io_memAXI_0_w_ready(io_memAXI_0_w_ready),
    .io_memAXI_0_w_valid(io_memAXI_0_w_valid),
    .io_memAXI_0_w_bits_data(io_memAXI_0_w_bits_data[0]),
    .io_memAXI_0_w_bits_strb(io_memAXI_0_w_bits_strb),
    .io_memAXI_0_w_bits_last(io_memAXI_0_w_bits_last),
    .io_memAXI_0_b_ready(io_memAXI_0_b_ready),
    .io_memAXI_0_b_valid(io_memAXI_0_b_valid),
    .io_memAXI_0_b_bits_resp(io_memAXI_0_b_bits_resp),
    .io_memAXI_0_b_bits_id(io_memAXI_0_b_bits_id),
    .io_memAXI_0_b_bits_user(io_memAXI_0_b_bits_user),
    .io_memAXI_0_ar_ready(io_memAXI_0_ar_ready),
    .io_memAXI_0_ar_valid(io_memAXI_0_ar_valid),
    .io_memAXI_0_ar_bits_addr(io_memAXI_0_ar_bits_addr),
    .io_memAXI_0_ar_bits_prot(io_memAXI_0_ar_bits_prot),
    .io_memAXI_0_ar_bits_id(io_memAXI_0_ar_bits_id),
    .io_memAXI_0_ar_bits_user(io_memAXI_0_ar_bits_user),
    .io_memAXI_0_ar_bits_len(io_memAXI_0_ar_bits_len),
    .io_memAXI_0_ar_bits_size(io_memAXI_0_ar_bits_size),
    .io_memAXI_0_ar_bits_burst(io_memAXI_0_ar_bits_burst),
    .io_memAXI_0_ar_bits_lock(io_memAXI_0_ar_bits_lock),
    .io_memAXI_0_ar_bits_cache(io_memAXI_0_ar_bits_cache),
    .io_memAXI_0_ar_bits_qos(io_memAXI_0_ar_bits_qos),
    .io_memAXI_0_r_ready(io_memAXI_0_r_ready),
    .io_memAXI_0_r_valid(io_memAXI_0_r_valid),
    .io_memAXI_0_r_bits_resp(io_memAXI_0_r_bits_resp),
    .io_memAXI_0_r_bits_data(io_memAXI_0_r_bits_data[0]),
    .io_memAXI_0_r_bits_last(io_memAXI_0_r_bits_last),
    .io_memAXI_0_r_bits_id(io_memAXI_0_r_bits_id),
    .io_memAXI_0_r_bits_user(io_memAXI_0_r_bits_user)
  );
endmodule
